class fifo_sequence extends uvm_sequence #(fifo_transaction);
  `uvm_object_utils(fifo_sequence) // Register the class with the factory

  // Declare handle to the transaction packet
  fifo_transaction tx;
  
  // Constructor 
  function new(string name="fifo_sequence");
    super.new(name);
  endfunction

  // virtual? 
  task body();
    if (starting_phase != null)
      starting_phase.raise_objection(this);

    // generate some transactions
    tx = fifo_transaction::type_id::create("tx");
    repeat(TX_COUNT_WR) begin
      start_item(tx);
      
      if (!tx.randomize())
        `uvm_error("RANDOMIZE", "Failed to randomize transaction")
      
      tx.wr_en = 1;
      tx.rd_en = 0;
      `uvm_info("GENERATE", tx.convert2string(), UVM_MEDIUM)
      finish_item(tx);
    end

    // generate some transactions
    repeat(TX_COUNT_RD) begin
      start_item(tx);
      
      tx.wr_en = 0;
      tx.rd_en = 1;
      `uvm_info("GENERATE", tx.convert2string(), UVM_MEDIUM)
      finish_item(tx);
    end



    if (starting_phase != null)
      starting_phase.drop_objection(this);
  endtask : body




endclass
