class scoreboard;
	
	// Instantiating the interface
	virtual Asynchronous_FIFO_bfm bfm;
	
	function new (virtual Asynchronous_FIFO_bfm b);
		bfm = b;
	endfunction
	
	task execute();
	
